
 /*
  Copyright 2013 Ray Salemi

  Licensed under the Apache License, Version 2.0 (the "License");
  you may not use this file except in compliance with the License.
  You may obtain a copy of the License at

  http://www.apache.org/licenses/LICENSE-2.0

  Unless required by applicable law or agreed to in writing, software
  distributed under the License is distributed on an "AS IS" BASIS,
  WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
  See the License for the specific language governing permissions and
  limitations under the License.
  */
 `timescale 1ns/1ps
package alu_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"

	typedef enum bit[2:0] {
		and_op  = 3'b000,
		or_op   = 3'b001,
		add_op  = 3'b100,
		sub_op  = 3'b101,
		rst_op  = 3'b110,
		no_op   = 3'b111 } operation_t;

	typedef struct packed {
		bit         signed  [31:0]  A;
		bit         signed  [31:0]  B;
		bit                 [3:0]   package_n;
		bit                         crc_ok;
		bit                 [3:0]   CRC;
		bit                 [3:0]   flags;
		bit                 [2:0]   crc_out;
		bit                         done;
		bit                 [5:0]   error;
		bit                         correct;
		bit                         sin;
		logic                       sout;
		operation_t                 op;
	} command_s;


`include "coverage.svh"
`include "base_tester.svh"
`include "random_tester.svh"
`include "corner_value_tester.svh"
`include "scoreboard.svh"
`include "driver.svh"
`include "command_monitor.svh"
`include "result_monitor.svh"
`include "env.svh"
`include "random_test.svh"
`include "corner_value_test.svh"


endpackage : alu_pkg
